ENTITY TESTBENCH2 IS
END TESTBENCH2;
ARCHITECTURE structure OF TESTBENCH2 IS
COMPONENT TESTER PORT(A:OUT BIT; C:IN BIT); END COMPONENT;
COMPONENT INVERTER2 PORT(A:IN BIT; C:OUT BIT); END COMPONENT;
SIGNAL A,C:BIT;
BEGIN
	tester1: TESTER PORT MAP (A,C);
	UUT: INVERTER2 PORT MAP (A,C);
END structure;