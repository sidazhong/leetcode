ENTITY testbench IS
END testbench;
ARCHITECTURE structure OF testbench IS
COMPONENT RS_tester PORT(R,S:OUT BIT; Q,QBAR:IN BIT); END COMPONENT;
COMPONENT RS PORT(R,s:IN BIT; Q,QBAR:OUT BIT); END COMPONENT;
SIGNAL R,S,Q,QBAR:BIT;
BEGIN
	tester: RS_tester PORT MAP (R,S,Q,QBAR);
	UUT: RS PORT MAP (R,S,Q,QBAR);
END structure;