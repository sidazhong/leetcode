ENTITY TESTBENCH4 IS
END TESTBENCH4;
ARCHITECTURE structure OF TESTBENCH4 IS
COMPONENT TESTER PORT(A:OUT BIT; C:IN BIT); END COMPONENT;
COMPONENT INVERTER4 PORT(A:IN BIT; C:OUT BIT); END COMPONENT;
SIGNAL A,C:BIT;
BEGIN
	tester1: TESTER PORT MAP (A,C);
	UUT: INVERTER4 PORT MAP (A,C);
END structure;