ENTITY EXOR IS
	PORT (a,b : IN BIT ; c : OUT BIT);
END EXOR;
ARCHITECTURE structure OF EXOR IS
COMPONENT ENOR1 PORT(a,b:IN BIT;c:OUT BIT); END COMPONENT;
COMPONENT ENOR2 PORT(a,b:IN BIT;c:OUT BIT); END COMPONENT;
COMPONENT ENOR3 PORT(a,b:IN BIT;c:OUT BIT); END COMPONENT;
COMPONENT ENOR4 PORT(a,b:IN BIT;c:OUT BIT); END COMPONENT;
COMPONENT ENOR5 PORT(a,b:IN BIT;c:OUT BIT); END COMPONENT;
SIGNAL e1,e2,e3,e4:BIT;
BEGIN
	ENOR1 PORT MAP (a,b,e1);
	ENOR2 PORT MAP (a,e1,e2);
	ENOR3 PORT MAP (b,e1,e3);
	ENOR4 PORT MAP (e2,e3,e4);
	ENOR5 PORT MAP (e4,e4,c);
END structure;