ENTITY INVERTER3 IS
	PORT (A : IN BIT ; C : OUT BIT);
END INVERTER3;
ARCHITECTURE structure OF INVERTER3 IS
COMPONENT ENOT_4 PORT(a:IN BIT;c:OUT BIT); END COMPONENT;
COMPONENT EAND_1 PORT(a,b:IN BIT;c:OUT BIT); END COMPONENT;
SIGNAL B:BIT;
BEGIN
	u1: ENOT_4 PORT MAP (A,B);
	u2: EAND_1 PORT MAP (A,B,C);
END structure;