ENTITY TESTBENCH3 IS
END TESTBENCH3;
ARCHITECTURE structure OF TESTBENCH3 IS
COMPONENT TESTER PORT(A:OUT BIT; C:IN BIT); END COMPONENT;
COMPONENT INVERTER3 PORT(A:IN BIT; C:OUT BIT); END COMPONENT;
SIGNAL A,C:BIT;
BEGIN
	tester1: TESTER PORT MAP (A,C);
	UUT: INVERTER3 PORT MAP (A,C);
END structure;