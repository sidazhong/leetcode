ENTITY TESTBENCH1 IS
END TESTBENCH1;
ARCHITECTURE structure OF TESTBENCH1 IS
COMPONENT TESTER PORT(A:OUT BIT; C:IN BIT); END COMPONENT;
COMPONENT INVERTER1 PORT(A:IN BIT; C:OUT BIT); END COMPONENT;
SIGNAL A,C:BIT;
BEGIN
	tester1: TESTER PORT MAP (A,C);
	UUT: INVERTER1 PORT MAP (A,C);
END structure;