ENTITY INVERTER4 IS
	PORT (A : IN BIT ; C : OUT BIT);
END INVERTER4;
ARCHITECTURE structure OF INVERTER4 IS
COMPONENT ENOT_4 PORT(a:IN BIT;c:OUT BIT); END COMPONENT;
COMPONENT EAND_3 PORT(a,b:IN BIT;c:OUT BIT); END COMPONENT;
SIGNAL B:BIT;
BEGIN
	u1: ENOT_4 PORT MAP (A,B);
	u2: EAND_3 PORT MAP (A,B,C);
END structure;