ENTITY RS IS
	PORT (R,S : IN BIT ; Q,QBAR : OUT BIT);
END RS;
ARCHITECTURE structure OF RS IS
COMPONENT ENOR1 PORT(a,b:IN BIT;c:OUT BIT); END COMPONENT;
COMPONENT ENOR2 PORT(a,b:IN BIT;c:OUT BIT); END COMPONENT;
BEGIN
	u1: ENOR1 PORT MAP (R,QBAR,Q);
	u2: ENOR2 PORT MAP (Q,S,QBAR);
END structure;